
module unsaved (
	vga_ball_0_clock_clk,
	audio_0_clk_clk,
	vga_ball_0_reset_reset,
	audio_0_reset_reset);	

	input		vga_ball_0_clock_clk;
	input		audio_0_clk_clk;
	input		vga_ball_0_reset_reset;
	input		audio_0_reset_reset;
endmodule
