`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Jakob Stiens
// 
// Create Date: 04/04/2022 04:37:56 PM
// Design Name: 
// Module Name: MegaShiftRegister
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module MegaShiftRegister #(parameter MSB = 9) (input clk, input logic enable, input logic direction, input logic [7:0] address,
                                            input logic [MSB:0] shift_in, output logic[MSB:0] outputData);

        wire[MSB:0] SRO1;
        wire[MSB:0] SRO2;
        wire[MSB:0] SRO3;
        wire[MSB:0] SRO4;
        wire[MSB:0] SRO5;
        wire[MSB:0] SRO6;
        wire[MSB:0] SRO7;
        wire[MSB:0] SRO8;
        wire[MSB:0] SRO9;
        wire[MSB:0] SRO10;
        wire[MSB:0] SRO11;
        wire[MSB:0] SRO12;
        wire[MSB:0] SRO13;
        wire[MSB:0] SRO14;
        wire[MSB:0] SRO15;
        wire[MSB:0] SRO16;
        wire[MSB:0] SRO17;
        wire[MSB:0] SRO18;
        wire[MSB:0] SRO19;
        wire[MSB:0] SRO20;
        wire[MSB:0] SRO21;
        wire[MSB:0] SRO22;
        wire[MSB:0] SRO23;
        wire[MSB:0] SRO24;
        wire[MSB:0] SRO25;
        wire[MSB:0] SRO26;
        wire[MSB:0] SRO27;
        wire[MSB:0] SRO28;
        wire[MSB:0] SRO29;
        wire[MSB:0] SRO30;
        wire[MSB:0] SRO31;
        wire[MSB:0] SRO32;
        wire[MSB:0] SRO33;
        wire[MSB:0] SRO34;
        wire[MSB:0] SRO35;
        wire[MSB:0] SRO36;
        wire[MSB:0] SRO37;
        wire[MSB:0] SRO38;
        wire[MSB:0] SRO39;
        wire[MSB:0] SRO40;
        wire[MSB:0] SRO41;
        wire[MSB:0] SRO42;
        wire[MSB:0] SRO43;
        wire[MSB:0] SRO44;
        wire[MSB:0] SRO45;
        wire[MSB:0] SRO46;
        wire[MSB:0] SRO47;
        wire[MSB:0] SRO48;
        wire[MSB:0] SRO49;
        wire[MSB:0] SRO50;
        wire[MSB:0] SRO51;
        wire[MSB:0] SRO52;
        wire[MSB:0] SRO53;
        wire[MSB:0] SRO54;
        wire[MSB:0] SRO55;
        wire[MSB:0] SRO56;
        wire[MSB:0] SRO57;
        wire[MSB:0] SRO58;
        wire[MSB:0] SRO59;
        wire[MSB:0] SRO60;
        wire[MSB:0] SRO61;
        wire[MSB:0] SRO62;
        wire[MSB:0] SRO63;
        wire[MSB:0] SRO64;
        wire[MSB:0] SRO65;
        wire[MSB:0] SRO66;
        wire[MSB:0] SRO67;
        wire[MSB:0] SRO68;
        wire[MSB:0] SRO69;
        wire[MSB:0] SRO70;
        wire[MSB:0] SRO71;
        wire[MSB:0] SRO72;
        wire[MSB:0] SRO73;
        wire[MSB:0] SRO74;
        wire[MSB:0] SRO75;
        wire[MSB:0] SRO76;
        wire[MSB:0] SRO77;
        wire[MSB:0] SRO78;
        wire[MSB:0] SRO79;
        wire[MSB:0] SRO80;
        wire[MSB:0] SRO81;
        wire[MSB:0] SRO82;
        wire[MSB:0] SRO83;
        wire[MSB:0] SRO84;
        wire[MSB:0] SRO85;
        wire[MSB:0] SRO86;
        wire[MSB:0] SRO87;
        wire[MSB:0] SRO88;
        wire[MSB:0] SRO89;
        wire[MSB:0] SRO90;
        wire[MSB:0] SRO91;
        wire[MSB:0] SRO92;
        wire[MSB:0] SRO93;
        wire[MSB:0] SRO94;
        wire[MSB:0] SRO95;
        wire[MSB:0] SRO96;
        wire[MSB:0] SRO97;
        wire[MSB:0] SRO98;
        wire[MSB:0] SRO99;
        wire[MSB:0] SRO100;
        wire[MSB:0] SRO101;
        wire[MSB:0] SRO102;
        wire[MSB:0] SRO103;
        wire[MSB:0] SRO104;
        wire[MSB:0] SRO105;
        wire[MSB:0] SRO106;
        wire[MSB:0] SRO107;
        wire[MSB:0] SRO108;
        wire[MSB:0] SRO109;
        wire[MSB:0] SRO110;
        wire[MSB:0] SRO111;
        wire[MSB:0] SRO112;
        wire[MSB:0] SRO113;
        wire[MSB:0] SRO114;
        wire[MSB:0] SRO115;
        wire[MSB:0] SRO116;
        wire[MSB:0] SRO117;
        wire[MSB:0] SRO118;
        wire[MSB:0] SRO119;
        wire[MSB:0] SRO120;
        wire[MSB:0] SRO121;
        wire[MSB:0] SRO122;
        wire[MSB:0] SRO123;
        wire[MSB:0] SRO124;
        wire[MSB:0] SRO125;
        wire[MSB:0] SRO126;
        wire[MSB:0] SRO127;
        wire[MSB:0] SRO128;
        wire[MSB:0] SRO129;
        wire[MSB:0] SRO130;
        wire[MSB:0] SRO131;
        wire[MSB:0] SRO132;
        wire[MSB:0] SRO133;
        wire[MSB:0] SRO134;
        wire[MSB:0] SRO135;
        wire[MSB:0] SRO136;
        wire[MSB:0] SRO137;
        wire[MSB:0] SRO138;
        wire[MSB:0] SRO139;
        wire[MSB:0] SRO140;
        wire[MSB:0] SRO141;
        wire[MSB:0] SRO142;
        wire[MSB:0] SRO143;
        wire[MSB:0] SRO144;
        wire[MSB:0] SRO145;
        wire[MSB:0] SRO146;
        wire[MSB:0] SRO147;
        wire[MSB:0] SRO148;
        wire[MSB:0] SRO149;
        wire[MSB:0] SRO150;
        wire[MSB:0] SRO151;
        wire[MSB:0] SRO152;
        wire[MSB:0] SRO153;
        wire[MSB:0] SRO154;
        wire[MSB:0] SRO155;
        wire[MSB:0] SRO156;
        wire[MSB:0] SRO157;
        wire[MSB:0] SRO158;
        wire[MSB:0] SRO159;
        wire[MSB:0] SRO160;
        wire[MSB:0] SRO161;
        wire[MSB:0] SRO162;
        wire[MSB:0] SRO163;
        wire[MSB:0] SRO164;
        wire[MSB:0] SRO165;
        wire[MSB:0] SRO166;
        wire[MSB:0] SRO167;
        wire[MSB:0] SRO168;
        wire[MSB:0] SRO169;
        wire[MSB:0] SRO170;
        wire[MSB:0] SRO171;
        wire[MSB:0] SRO172;
        wire[MSB:0] SRO173;
        wire[MSB:0] SRO174;
        wire[MSB:0] SRO175;
        wire[MSB:0] SRO176;
        wire[MSB:0] SRO177;
        wire[MSB:0] SRO178;
        wire[MSB:0] SRO179;
        wire[MSB:0] SRO180;
        wire[MSB:0] SRO181;
        wire[MSB:0] SRO182;
        wire[MSB:0] SRO183;
        wire[MSB:0] SRO184;
        wire[MSB:0] SRO185;
        wire[MSB:0] SRO186;
        wire[MSB:0] SRO187;
        wire[MSB:0] SRO188;
        wire[MSB:0] SRO189;
        wire[MSB:0] SRO190;
        wire[MSB:0] SRO191;
        wire[MSB:0] SRO192;
        wire[MSB:0] SRO193;
        wire[MSB:0] SRO194;
        wire[MSB:0] SRO195;
        wire[MSB:0] SRO196;
        wire[MSB:0] SRO197;
        wire[MSB:0] SRO198;
        wire[MSB:0] SRO199;
        wire[MSB:0] SRO200;
        wire[MSB:0] SRO201;
        wire[MSB:0] SRO202;
        wire[MSB:0] SRO203;
        wire[MSB:0] SRO204;
        wire[MSB:0] SRO205;
        wire[MSB:0] SRO206;
        wire[MSB:0] SRO207;
        wire[MSB:0] SRO208;
        wire[MSB:0] SRO209;
        wire[MSB:0] SRO210;
        wire[MSB:0] SRO211;
        wire[MSB:0] SRO212;
        wire[MSB:0] SRO213;
        wire[MSB:0] SRO214;
        wire[MSB:0] SRO215;
        wire[MSB:0] SRO216;
        wire[MSB:0] SRO217;
        wire[MSB:0] SRO218;
        wire[MSB:0] SRO219;
        wire[MSB:0] SRO220;
        wire[MSB:0] SRO221;
        wire[MSB:0] SRO222;
        wire[MSB:0] SRO223;
        wire[MSB:0] SRO224;
        wire[MSB:0] SRO225;
        wire[MSB:0] SRO226;
        wire[MSB:0] SRO227;
        wire[MSB:0] SRO228;
        wire[MSB:0] SRO229;
        wire[MSB:0] SRO230;
        wire[MSB:0] SRO231;
        wire[MSB:0] SRO232;
        wire[MSB:0] SRO233;
        wire[MSB:0] SRO234;
        wire[MSB:0] SRO235;
        wire[MSB:0] SRO236;
        wire[MSB:0] SRO237;
        wire[MSB:0] SRO238;
        wire[MSB:0] SRO239;
        wire[MSB:0] SRO240;

        shift_register SR1(.clk(clk), .enable(enable), .direction(direction), .reset(reset), 
                                            .data(shift_in), .outputData(SRO1));
        shift_register SR2(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO1), .outputData(SRO2));
        shift_register SR3(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO2), .outputData(SRO3));
        shift_register SR4(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO3), .outputData(SRO4));
        shift_register SR5(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO4), .outputData(SRO5));
        shift_register SR6(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO5), .outputData(SRO6));
        shift_register SR7(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO6), .outputData(SRO7));
        shift_register SR8(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO7), .outputData(SRO8));
        shift_register SR9(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO8), .outputData(SRO9));
        shift_register SR10(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO9), .outputData(SRO10));
        shift_register SR11(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO10), .outputData(SRO11));
        shift_register SR12(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO11), .outputData(SRO12));
        shift_register SR13(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO12), .outputData(SRO13));
        shift_register SR14(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO13), .outputData(SRO14));
        shift_register SR15(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO14), .outputData(SRO15));
        shift_register SR16(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO15), .outputData(SRO16));
        shift_register SR17(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO16), .outputData(SRO17));
        shift_register SR18(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO17), .outputData(SRO18));
        shift_register SR19(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO18), .outputData(SRO19));
        shift_register SR20(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO19), .outputData(SRO20));
        shift_register SR21(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO20), .outputData(SRO21));
        shift_register SR22(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO21), .outputData(SRO22));
        shift_register SR23(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO22), .outputData(SRO23));
        shift_register SR24(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO23), .outputData(SRO24));
        shift_register SR25(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO24), .outputData(SRO25));
        shift_register SR26(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO25), .outputData(SRO26));
        shift_register SR27(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO26), .outputData(SRO27));
        shift_register SR28(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO27), .outputData(SRO28));
        shift_register SR29(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO28), .outputData(SRO29));
        shift_register SR30(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO29), .outputData(SRO30));
        shift_register SR31(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO30), .outputData(SRO31));
        shift_register SR32(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO31), .outputData(SRO32));
        shift_register SR33(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO32), .outputData(SRO33));
        shift_register SR34(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO33), .outputData(SRO34));
        shift_register SR35(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO34), .outputData(SRO35));
        shift_register SR36(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO35), .outputData(SRO36));
        shift_register SR37(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO36), .outputData(SRO37));
        shift_register SR38(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO37), .outputData(SRO38));
        shift_register SR39(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO38), .outputData(SRO39));
        shift_register SR40(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO39), .outputData(SRO40));
        shift_register SR41(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO40), .outputData(SRO41));
        shift_register SR42(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO41), .outputData(SRO42));
        shift_register SR43(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO42), .outputData(SRO43));
        shift_register SR44(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO43), .outputData(SRO44));
        shift_register SR45(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO44), .outputData(SRO45));
        shift_register SR46(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO45), .outputData(SRO46));
        shift_register SR47(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO46), .outputData(SRO47));
        shift_register SR48(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO47), .outputData(SRO48));
        shift_register SR49(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO48), .outputData(SRO49));
        shift_register SR50(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO49), .outputData(SRO50));
        shift_register SR51(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO50), .outputData(SRO51));
        shift_register SR52(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO51), .outputData(SRO52));
        shift_register SR53(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO52), .outputData(SRO53));
        shift_register SR54(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO53), .outputData(SRO54));
        shift_register SR55(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO54), .outputData(SRO55));
        shift_register SR56(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO55), .outputData(SRO56));
        shift_register SR57(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO56), .outputData(SRO57));
        shift_register SR58(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO57), .outputData(SRO58));
        shift_register SR59(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO58), .outputData(SRO59));
        shift_register SR60(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO59), .outputData(SRO60));
        shift_register SR61(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO60), .outputData(SRO61));
        shift_register SR62(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO61), .outputData(SRO62));
        shift_register SR63(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO62), .outputData(SRO63));
        shift_register SR64(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO63), .outputData(SRO64));
        shift_register SR65(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO64), .outputData(SRO65));
        shift_register SR66(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO65), .outputData(SRO66));
        shift_register SR67(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO66), .outputData(SRO67));
        shift_register SR68(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO67), .outputData(SRO68));
        shift_register SR69(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO68), .outputData(SRO69));
        shift_register SR70(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO69), .outputData(SRO70));
        shift_register SR71(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO70), .outputData(SRO71));
        shift_register SR72(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO71), .outputData(SRO72));
        shift_register SR73(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO72), .outputData(SRO73));
        shift_register SR74(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO73), .outputData(SRO74));
        shift_register SR75(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO74), .outputData(SRO75));
        shift_register SR76(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO75), .outputData(SRO76));
        shift_register SR77(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO76), .outputData(SRO77));
        shift_register SR78(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO77), .outputData(SRO78));
        shift_register SR79(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO78), .outputData(SRO79));
        shift_register SR80(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO79), .outputData(SRO80));
        shift_register SR81(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO80), .outputData(SRO81));
        shift_register SR82(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO81), .outputData(SRO82));
        shift_register SR83(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO82), .outputData(SRO83));
        shift_register SR84(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO83), .outputData(SRO84));
        shift_register SR85(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO84), .outputData(SRO85));
        shift_register SR86(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO85), .outputData(SRO86));
        shift_register SR87(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO86), .outputData(SRO87));
        shift_register SR88(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO87), .outputData(SRO88));
        shift_register SR89(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO88), .outputData(SRO89));
        shift_register SR90(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO89), .outputData(SRO90));
        shift_register SR91(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO90), .outputData(SRO91));
        shift_register SR92(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO91), .outputData(SRO92));
        shift_register SR93(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO92), .outputData(SRO93));
        shift_register SR94(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO93), .outputData(SRO94));
        shift_register SR95(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO94), .outputData(SRO95));
        shift_register SR96(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO95), .outputData(SRO96));
        shift_register SR97(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO96), .outputData(SRO97));
        shift_register SR98(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO97), .outputData(SRO98));
        shift_register SR99(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO98), .outputData(SRO99));
        shift_register SR100(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO99), .outputData(SRO100));
        shift_register SR101(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO100), .outputData(SRO101));
        shift_register SR102(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO101), .outputData(SRO102));
        shift_register SR103(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO102), .outputData(SRO103));
        shift_register SR104(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO103), .outputData(SRO104));
        shift_register SR105(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO104), .outputData(SRO105));
        shift_register SR106(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO105), .outputData(SRO106));
        shift_register SR107(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO106), .outputData(SRO107));
        shift_register SR108(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO107), .outputData(SRO108));
        shift_register SR109(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO108), .outputData(SRO109));
        shift_register SR110(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO109), .outputData(SRO110));
        shift_register SR111(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO110), .outputData(SRO111));
        shift_register SR112(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO111), .outputData(SRO112));
        shift_register SR113(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO112), .outputData(SRO113));
        shift_register SR114(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO113), .outputData(SRO114));
        shift_register SR115(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO114), .outputData(SRO115));
        shift_register SR116(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO115), .outputData(SRO116));
        shift_register SR117(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO116), .outputData(SRO117));
        shift_register SR118(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO117), .outputData(SRO118));
        shift_register SR119(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO118), .outputData(SRO119));
        shift_register SR120(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO119), .outputData(SRO120));
        shift_register SR121(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO120), .outputData(SRO121));
        shift_register SR122(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO121), .outputData(SRO122));
        shift_register SR123(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO122), .outputData(SRO123));
        shift_register SR124(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO123), .outputData(SRO124));
        shift_register SR125(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO124), .outputData(SRO125));
        shift_register SR126(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO125), .outputData(SRO126));
        shift_register SR127(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO126), .outputData(SRO127));
        shift_register SR128(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO127), .outputData(SRO128));
        shift_register SR129(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO128), .outputData(SRO129));
        shift_register SR130(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO129), .outputData(SRO130));
        shift_register SR131(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO130), .outputData(SRO131));
        shift_register SR132(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO131), .outputData(SRO132));
        shift_register SR133(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO132), .outputData(SRO133));
        shift_register SR134(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO133), .outputData(SRO134));
        shift_register SR135(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO134), .outputData(SRO135));
        shift_register SR136(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO135), .outputData(SRO136));
        shift_register SR137(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO136), .outputData(SRO137));
        shift_register SR138(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO137), .outputData(SRO138));
        shift_register SR139(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO138), .outputData(SRO139));
        shift_register SR140(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO139), .outputData(SRO140));
        shift_register SR141(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO140), .outputData(SRO141));
        shift_register SR142(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO141), .outputData(SRO142));
        shift_register SR143(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO142), .outputData(SRO143));
        shift_register SR144(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO143), .outputData(SRO144));
        shift_register SR145(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO144), .outputData(SRO145));
        shift_register SR146(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO145), .outputData(SRO146));
        shift_register SR147(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO146), .outputData(SRO147));
        shift_register SR148(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO147), .outputData(SRO148));
        shift_register SR149(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO148), .outputData(SRO149));
        shift_register SR150(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO149), .outputData(SRO150));
        shift_register SR151(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO150), .outputData(SRO151));
        shift_register SR152(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO151), .outputData(SRO152));
        shift_register SR153(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO152), .outputData(SRO153));
        shift_register SR154(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO153), .outputData(SRO154));
        shift_register SR155(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO154), .outputData(SRO155));
        shift_register SR156(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO155), .outputData(SRO156));
        shift_register SR157(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO156), .outputData(SRO157));
        shift_register SR158(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO157), .outputData(SRO158));
        shift_register SR159(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO158), .outputData(SRO159));
        shift_register SR160(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO159), .outputData(SRO160));
        shift_register SR161(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO160), .outputData(SRO161));
        shift_register SR162(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO161), .outputData(SRO162));
        shift_register SR163(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO162), .outputData(SRO163));
        shift_register SR164(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO163), .outputData(SRO164));
        shift_register SR165(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO164), .outputData(SRO165));
        shift_register SR166(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO165), .outputData(SRO166));
        shift_register SR167(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO166), .outputData(SRO167));
        shift_register SR168(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO167), .outputData(SRO168));
        shift_register SR169(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO168), .outputData(SRO169));
        shift_register SR170(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO169), .outputData(SRO170));
        shift_register SR171(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO170), .outputData(SRO171));
        shift_register SR172(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO171), .outputData(SRO172));
        shift_register SR173(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO172), .outputData(SRO173));
        shift_register SR174(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO173), .outputData(SRO174));
        shift_register SR175(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO174), .outputData(SRO175));
        shift_register SR176(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO175), .outputData(SRO176));
        shift_register SR177(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO176), .outputData(SRO177));
        shift_register SR178(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO177), .outputData(SRO178));
        shift_register SR179(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO178), .outputData(SRO179));
        shift_register SR180(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO179), .outputData(SRO180));
        shift_register SR181(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO180), .outputData(SRO181));
        shift_register SR182(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO181), .outputData(SRO182));
        shift_register SR183(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO182), .outputData(SRO183));
        shift_register SR184(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO183), .outputData(SRO184));
        shift_register SR185(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO184), .outputData(SRO185));
        shift_register SR186(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO185), .outputData(SRO186));
        shift_register SR187(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO186), .outputData(SRO187));
        shift_register SR188(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO187), .outputData(SRO188));
        shift_register SR189(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO188), .outputData(SRO189));
        shift_register SR190(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO189), .outputData(SRO190));
        shift_register SR191(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO190), .outputData(SRO191));
        shift_register SR192(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO191), .outputData(SRO192));
        shift_register SR193(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO192), .outputData(SRO193));
        shift_register SR194(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO193), .outputData(SRO194));
        shift_register SR195(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO194), .outputData(SRO195));
        shift_register SR196(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO195), .outputData(SRO196));
        shift_register SR197(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO196), .outputData(SRO197));
        shift_register SR198(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO197), .outputData(SRO198));
        shift_register SR199(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO198), .outputData(SRO199));
        shift_register SR200(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO199), .outputData(SRO200));
        shift_register SR201(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO200), .outputData(SRO201));
        shift_register SR202(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO201), .outputData(SRO202));
        shift_register SR203(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO202), .outputData(SRO203));
        shift_register SR204(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO203), .outputData(SRO204));
        shift_register SR205(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO204), .outputData(SRO205));
        shift_register SR206(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO205), .outputData(SRO206));
        shift_register SR207(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO206), .outputData(SRO207));
        shift_register SR208(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO207), .outputData(SRO208));
        shift_register SR209(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO208), .outputData(SRO209));
        shift_register SR210(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO209), .outputData(SRO210));
        shift_register SR211(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO210), .outputData(SRO211));
        shift_register SR212(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO211), .outputData(SRO212));
        shift_register SR213(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO212), .outputData(SRO213));
        shift_register SR214(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO213), .outputData(SRO214));
        shift_register SR215(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO214), .outputData(SRO215));
        shift_register SR216(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO215), .outputData(SRO216));
        shift_register SR217(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO216), .outputData(SRO217));
        shift_register SR218(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO217), .outputData(SRO218));
        shift_register SR219(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO218), .outputData(SRO219));
        shift_register SR220(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO219), .outputData(SRO220));
        shift_register SR221(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO220), .outputData(SRO221));
        shift_register SR222(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO221), .outputData(SRO222));
        shift_register SR223(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO222), .outputData(SRO223));
        shift_register SR224(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO223), .outputData(SRO224));
        shift_register SR225(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO224), .outputData(SRO225));
        shift_register SR226(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO225), .outputData(SRO226));
        shift_register SR227(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO226), .outputData(SRO227));
        shift_register SR228(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO227), .outputData(SRO228));
        shift_register SR229(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO228), .outputData(SRO229));
        shift_register SR230(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO229), .outputData(SRO230));
        shift_register SR231(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO230), .outputData(SRO231));
        shift_register SR232(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO231), .outputData(SRO232));
        shift_register SR233(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO232), .outputData(SRO233));
        shift_register SR234(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO233), .outputData(SRO234));
        shift_register SR235(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO234), .outputData(SRO235));
        shift_register SR236(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO235), .outputData(SRO236));
        shift_register SR237(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO236), .outputData(SRO237));
        shift_register SR238(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO237), .outputData(SRO238));
        shift_register SR239(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO238), .outputData(SRO239));
        shift_register SR240(.clk(clk), .enable(enable), .direction(direction), .reset(reset), .data(SRO239), .outputData(SRO240));


        logic [MSB:0] outputDataStore;
        
        assign outputData = outputDataStore; 
        
        always @(posedge clk) begin
            case (address)
            
                0 :  outputDataStore <= SRO1[MSB:0];
                1 :  outputDataStore <= SRO2[MSB:0];
                2 :  outputDataStore <= SRO3[MSB:0];
                3 :  outputDataStore <= SRO4[MSB:0];
                4 :  outputDataStore <= SRO5[MSB:0];
                5 :  outputDataStore <= SRO6[MSB:0];
                6 :  outputDataStore <= SRO7[MSB:0];
                7 :  outputDataStore <= SRO8[MSB:0];
                8 :  outputDataStore <= SRO9[MSB:0];
                9 :  outputDataStore <= SRO10[MSB:0];
                10 :  outputDataStore <= SRO11[MSB:0];
                11 :  outputDataStore <= SRO12[MSB:0];
                12 :  outputDataStore <= SRO13[MSB:0];
                13 :  outputDataStore <= SRO14[MSB:0];
                14 :  outputDataStore <= SRO15[MSB:0];
                15 :  outputDataStore <= SRO16[MSB:0];
                16 :  outputDataStore <= SRO17[MSB:0];
                17 :  outputDataStore <= SRO18[MSB:0];
                18 :  outputDataStore <= SRO19[MSB:0];
                19 :  outputDataStore <= SRO20[MSB:0];
                20 :  outputDataStore <= SRO21[MSB:0];
                21 :  outputDataStore <= SRO22[MSB:0];
                22 :  outputDataStore <= SRO23[MSB:0];
                23 :  outputDataStore <= SRO24[MSB:0];
                24 :  outputDataStore <= SRO25[MSB:0];
                25 :  outputDataStore <= SRO26[MSB:0];
                26 :  outputDataStore <= SRO27[MSB:0];
                27 :  outputDataStore <= SRO28[MSB:0];
                28 :  outputDataStore <= SRO29[MSB:0];
                29 :  outputDataStore <= SRO30[MSB:0];
                30 :  outputDataStore <= SRO31[MSB:0];
                31 :  outputDataStore <= SRO32[MSB:0];
                32 :  outputDataStore <= SRO33[MSB:0];
                33 :  outputDataStore <= SRO34[MSB:0];
                34 :  outputDataStore <= SRO35[MSB:0];
                35 :  outputDataStore <= SRO36[MSB:0];
                36 :  outputDataStore <= SRO37[MSB:0];
                37 :  outputDataStore <= SRO38[MSB:0];
                38 :  outputDataStore <= SRO39[MSB:0];
                39 :  outputDataStore <= SRO40[MSB:0];
                40 :  outputDataStore <= SRO41[MSB:0];
                41 :  outputDataStore <= SRO42[MSB:0];
                42 :  outputDataStore <= SRO43[MSB:0];
                43 :  outputDataStore <= SRO44[MSB:0];
                44 :  outputDataStore <= SRO45[MSB:0];
                45 :  outputDataStore <= SRO46[MSB:0];
                46 :  outputDataStore <= SRO47[MSB:0];
                47 :  outputDataStore <= SRO48[MSB:0];
                48 :  outputDataStore <= SRO49[MSB:0];
                49 :  outputDataStore <= SRO50[MSB:0];
                50 :  outputDataStore <= SRO51[MSB:0];
                51 :  outputDataStore <= SRO52[MSB:0];
                52 :  outputDataStore <= SRO53[MSB:0];
                53 :  outputDataStore <= SRO54[MSB:0];
                54 :  outputDataStore <= SRO55[MSB:0];
                55 :  outputDataStore <= SRO56[MSB:0];
                56 :  outputDataStore <= SRO57[MSB:0];
                57 :  outputDataStore <= SRO58[MSB:0];
                58 :  outputDataStore <= SRO59[MSB:0];
                59 :  outputDataStore <= SRO60[MSB:0];
                60 :  outputDataStore <= SRO61[MSB:0];
                61 :  outputDataStore <= SRO62[MSB:0];
                62 :  outputDataStore <= SRO63[MSB:0];
                63 :  outputDataStore <= SRO64[MSB:0];
                64 :  outputDataStore <= SRO65[MSB:0];
                65 :  outputDataStore <= SRO66[MSB:0];
                66 :  outputDataStore <= SRO67[MSB:0];
                67 :  outputDataStore <= SRO68[MSB:0];
                68 :  outputDataStore <= SRO69[MSB:0];
                69 :  outputDataStore <= SRO70[MSB:0];
                70 :  outputDataStore <= SRO71[MSB:0];
                71 :  outputDataStore <= SRO72[MSB:0];
                72 :  outputDataStore <= SRO73[MSB:0];
                73 :  outputDataStore <= SRO74[MSB:0];
                74 :  outputDataStore <= SRO75[MSB:0];
                75 :  outputDataStore <= SRO76[MSB:0];
                76 :  outputDataStore <= SRO77[MSB:0];
                77 :  outputDataStore <= SRO78[MSB:0];
                78 :  outputDataStore <= SRO79[MSB:0];
                79 :  outputDataStore <= SRO80[MSB:0];
                80 :  outputDataStore <= SRO81[MSB:0];
                81 :  outputDataStore <= SRO82[MSB:0];
                82 :  outputDataStore <= SRO83[MSB:0];
                83 :  outputDataStore <= SRO84[MSB:0];
                84 :  outputDataStore <= SRO85[MSB:0];
                85 :  outputDataStore <= SRO86[MSB:0];
                86 :  outputDataStore <= SRO87[MSB:0];
                87 :  outputDataStore <= SRO88[MSB:0];
                88 :  outputDataStore <= SRO89[MSB:0];
                89 :  outputDataStore <= SRO90[MSB:0];
                90 :  outputDataStore <= SRO91[MSB:0];
                91 :  outputDataStore <= SRO92[MSB:0];
                92 :  outputDataStore <= SRO93[MSB:0];
                93 :  outputDataStore <= SRO94[MSB:0];
                94 :  outputDataStore <= SRO95[MSB:0];
                95 :  outputDataStore <= SRO96[MSB:0];
                96 :  outputDataStore <= SRO97[MSB:0];
                97 :  outputDataStore <= SRO98[MSB:0];
                98 :  outputDataStore <= SRO99[MSB:0];
                99 :  outputDataStore <= SRO100[MSB:0];
                100 :  outputDataStore <= SRO101[MSB:0];
                101 :  outputDataStore <= SRO102[MSB:0];
                102 :  outputDataStore <= SRO103[MSB:0];
                103 :  outputDataStore <= SRO104[MSB:0];
                104 :  outputDataStore <= SRO105[MSB:0];
                105 :  outputDataStore <= SRO106[MSB:0];
                106 :  outputDataStore <= SRO107[MSB:0];
                107 :  outputDataStore <= SRO108[MSB:0];
                108 :  outputDataStore <= SRO109[MSB:0];
                109 :  outputDataStore <= SRO110[MSB:0];
                110 :  outputDataStore <= SRO111[MSB:0];
                111 :  outputDataStore <= SRO112[MSB:0];
                112 :  outputDataStore <= SRO113[MSB:0];
                113 :  outputDataStore <= SRO114[MSB:0];
                114 :  outputDataStore <= SRO115[MSB:0];
                115 :  outputDataStore <= SRO116[MSB:0];
                116 :  outputDataStore <= SRO117[MSB:0];
                117 :  outputDataStore <= SRO118[MSB:0];
                118 :  outputDataStore <= SRO119[MSB:0];
                119 :  outputDataStore <= SRO120[MSB:0];
                120 :  outputDataStore <= SRO121[MSB:0];
                121 :  outputDataStore <= SRO122[MSB:0];
                122 :  outputDataStore <= SRO123[MSB:0];
                123 :  outputDataStore <= SRO124[MSB:0];
                124 :  outputDataStore <= SRO125[MSB:0];
                125 :  outputDataStore <= SRO126[MSB:0];
                126 :  outputDataStore <= SRO127[MSB:0];
                127 :  outputDataStore <= SRO128[MSB:0];
                128 :  outputDataStore <= SRO129[MSB:0];
                129 :  outputDataStore <= SRO130[MSB:0];
                130 :  outputDataStore <= SRO131[MSB:0];
                131 :  outputDataStore <= SRO132[MSB:0];
                132 :  outputDataStore <= SRO133[MSB:0];
                133 :  outputDataStore <= SRO134[MSB:0];
                134 :  outputDataStore <= SRO135[MSB:0];
                135 :  outputDataStore <= SRO136[MSB:0];
                136 :  outputDataStore <= SRO137[MSB:0];
                137 :  outputDataStore <= SRO138[MSB:0];
                138 :  outputDataStore <= SRO139[MSB:0];
                139 :  outputDataStore <= SRO140[MSB:0];
                140 :  outputDataStore <= SRO141[MSB:0];
                141 :  outputDataStore <= SRO142[MSB:0];
                142 :  outputDataStore <= SRO143[MSB:0];
                143 :  outputDataStore <= SRO144[MSB:0];
                144 :  outputDataStore <= SRO145[MSB:0];
                145 :  outputDataStore <= SRO146[MSB:0];
                146 :  outputDataStore <= SRO147[MSB:0];
                147 :  outputDataStore <= SRO148[MSB:0];
                148 :  outputDataStore <= SRO149[MSB:0];
                149 :  outputDataStore <= SRO150[MSB:0];
                150 :  outputDataStore <= SRO151[MSB:0];
                151 :  outputDataStore <= SRO152[MSB:0];
                152 :  outputDataStore <= SRO153[MSB:0];
                153 :  outputDataStore <= SRO154[MSB:0];
                154 :  outputDataStore <= SRO155[MSB:0];
                155 :  outputDataStore <= SRO156[MSB:0];
                156 :  outputDataStore <= SRO157[MSB:0];
                157 :  outputDataStore <= SRO158[MSB:0];
                158 :  outputDataStore <= SRO159[MSB:0];
                159 :  outputDataStore <= SRO160[MSB:0];
                160 :  outputDataStore <= SRO161[MSB:0];
                161 :  outputDataStore <= SRO162[MSB:0];
                162 :  outputDataStore <= SRO163[MSB:0];
                163 :  outputDataStore <= SRO164[MSB:0];
                164 :  outputDataStore <= SRO165[MSB:0];
                165 :  outputDataStore <= SRO166[MSB:0];
                166 :  outputDataStore <= SRO167[MSB:0];
                167 :  outputDataStore <= SRO168[MSB:0];
                168 :  outputDataStore <= SRO169[MSB:0];
                169 :  outputDataStore <= SRO170[MSB:0];
                170 :  outputDataStore <= SRO171[MSB:0];
                171 :  outputDataStore <= SRO172[MSB:0];
                172 :  outputDataStore <= SRO173[MSB:0];
                173 :  outputDataStore <= SRO174[MSB:0];
                174 :  outputDataStore <= SRO175[MSB:0];
                175 :  outputDataStore <= SRO176[MSB:0];
                176 :  outputDataStore <= SRO177[MSB:0];
                177 :  outputDataStore <= SRO178[MSB:0];
                178 :  outputDataStore <= SRO179[MSB:0];
                179 :  outputDataStore <= SRO180[MSB:0];
                180 :  outputDataStore <= SRO181[MSB:0];
                181 :  outputDataStore <= SRO182[MSB:0];
                182 :  outputDataStore <= SRO183[MSB:0];
                183 :  outputDataStore <= SRO184[MSB:0];
                184 :  outputDataStore <= SRO185[MSB:0];
                185 :  outputDataStore <= SRO186[MSB:0];
                186 :  outputDataStore <= SRO187[MSB:0];
                187 :  outputDataStore <= SRO188[MSB:0];
                188 :  outputDataStore <= SRO189[MSB:0];
                189 :  outputDataStore <= SRO190[MSB:0];
                190 :  outputDataStore <= SRO191[MSB:0];
                191 :  outputDataStore <= SRO192[MSB:0];
                192 :  outputDataStore <= SRO193[MSB:0];
                193 :  outputDataStore <= SRO194[MSB:0];
                194 :  outputDataStore <= SRO195[MSB:0];
                195 :  outputDataStore <= SRO196[MSB:0];
                196 :  outputDataStore <= SRO197[MSB:0];
                197 :  outputDataStore <= SRO198[MSB:0];
                198 :  outputDataStore <= SRO199[MSB:0];
                199 :  outputDataStore <= SRO200[MSB:0];
                200 :  outputDataStore <= SRO201[MSB:0];
                201 :  outputDataStore <= SRO202[MSB:0];
                202 :  outputDataStore <= SRO203[MSB:0];
                203 :  outputDataStore <= SRO204[MSB:0];
                204 :  outputDataStore <= SRO205[MSB:0];
                205 :  outputDataStore <= SRO206[MSB:0];
                206 :  outputDataStore <= SRO207[MSB:0];
                207 :  outputDataStore <= SRO208[MSB:0];
                208 :  outputDataStore <= SRO209[MSB:0];
                209 :  outputDataStore <= SRO210[MSB:0];
                210 :  outputDataStore <= SRO211[MSB:0];
                211 :  outputDataStore <= SRO212[MSB:0];
                212 :  outputDataStore <= SRO213[MSB:0];
                213 :  outputDataStore <= SRO214[MSB:0];
                214 :  outputDataStore <= SRO215[MSB:0];
                215 :  outputDataStore <= SRO216[MSB:0];
                216 :  outputDataStore <= SRO217[MSB:0];
                217 :  outputDataStore <= SRO218[MSB:0];
                218 :  outputDataStore <= SRO219[MSB:0];
                219 :  outputDataStore <= SRO220[MSB:0];
                220 :  outputDataStore <= SRO221[MSB:0];
                221 :  outputDataStore <= SRO222[MSB:0];
                222 :  outputDataStore <= SRO223[MSB:0];
                223 :  outputDataStore <= SRO224[MSB:0];
                224 :  outputDataStore <= SRO225[MSB:0];
                225 :  outputDataStore <= SRO226[MSB:0];
                226 :  outputDataStore <= SRO227[MSB:0];
                227 :  outputDataStore <= SRO228[MSB:0];
                228 :  outputDataStore <= SRO229[MSB:0];
                229 :  outputDataStore <= SRO230[MSB:0];
                230 :  outputDataStore <= SRO231[MSB:0];
                231 :  outputDataStore <= SRO232[MSB:0];
                232 :  outputDataStore <= SRO233[MSB:0];
                233 :  outputDataStore <= SRO234[MSB:0];
                234 :  outputDataStore <= SRO235[MSB:0];
                235 :  outputDataStore <= SRO236[MSB:0];
                236 :  outputDataStore <= SRO237[MSB:0];
                237 :  outputDataStore <= SRO238[MSB:0];
                238 :  outputDataStore <= SRO239[MSB:0];
                239 :  outputDataStore <= SRO240[MSB:0];

                default : outputDataStore <= 5;
                
            endcase
        end 
        
        
        
                                               
endmodule
