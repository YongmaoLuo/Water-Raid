/*
 * Avalon memory-mapped peripheral that generates VGA
 *
 * Stephen A. Edwards
 * Columbia University
 */

module vga(	input logic        clk,
	        input logic 	   reset,
		input logic [15:0]  writedata,
		input logic 	   write,
		input 		   chipselect,
		input logic [5:0]  address,

		output logic [3:0] VGA_R, VGA_G, VGA_B,
		output logic 	   VGA_CLK, VGA_HS, VGA_VS,
		                   VGA_BLANK_n,
		output logic 	   VGA_SYNC_n);f

   logic [10:0]	   hcount;
   logic [9:0]     vcount;
   
   logic [9:0]	   boundary_1;
   logic [9:0]	   boundary_2;
   logic [9:0]	   boundary_3;
   logic [9:0]	   boundary_4;

   // last bit of y positions indicates whether sprite is onscreen

   logic [9:0]	   plane_x;
   logic [9:0]	   plane_y;

   logic [9:0]	   enemy_1_x;
   logic [9:0]	   enemy_1_y;

   logic [9:0]	   enemy_2_x;
   logic [9:0]	   enemy_2_y;

   logic [9:0]	   enemy_3_x;
   logic [9:0]	   enemy_3_y;

   logic [9:0]	   enemy_4_x;
   logic [9:0]	   enemy_4_y;

   logic [9:0]	   enemy_5_x;
   logic [9:0]	   enemy_5_y;

   logic [9:0]	   enemy_6_x;
   logic [9:0]	   enemy_6_y;

   logic [9:0]	   enemy_7_x;
   logic [9:0]	   enemy_7_y;

   logic [9:0]	   enemy_8_x;
   logic [9:0]	   enemy_8_y;

   logic [9:0]	   bullet_x;
   logic [9:0]	   bullet_y;

   logic [9:0]	   explosion_x;
   logic [9:0]	   explosion_y;

   logic [3:0]	   score_digit_1;
   logic [3:0]	   score_digit_2;
   logic [3:0]	   score_digit_3;
   logic [3:0]	   score_digit_4;
   logic [3:0]	   score_digit_5;

   logic	   isMusic;
   logic [1:0]	   whichClip;

   logic [7:0] 	   background_r, background_g, background_b;
	
   vga_counters counters(.clk50(clk), .*);

   always_ff @(posedge clk)
     if (reset) begin
	background_r <= 8'h0;
	background_g <= 8'h0;
	background_b <= 8'h80;
     end else if (chipselect && write)
       case (address)
	 6'h0 : background_r <= writedata[3:0];
	 6'h1 : background_g <= writedata[3:0];
	 6'h2 : background_b <= writedata[3:0]; 
	 6'h3 : boundary_1 <= writedata[9:0];
	 6'h4 : boundary_2 <= writedata[9:0];
	 6'h5 : boundary_3 <= writedata[9:0];
	 6'h6 : boundary_4 <= writedata[9:0];
	 6'h7 : plane_x <= writedata[9:0]; 
	 6'h8 : plane_y <= writedata[9:0];
   	 6'h9 : enemy_1_x <= writedata[9:0];
   	 6'h10 : enemy_1_y <= writedata[9:0];
         6'h12 : enemy_2_x <= writedata[9:0];
         6'h13 : enemy_2_y <= writedata[9:0];
         6'h14 : enemy_3_x <= writedata[9:0];
         6'h15 : enemy_3_y <= writedata[9:0];
         6'h16 : enemy_4_x <= writedata[9:0];
         6'h17 : enemy_4_y <= writedata[9:0];
         6'h18 : enemy_5_x <= writedata[9:0];
         6'h19 : enemy_5_y <= writedata[9:0];
         6'h20 : enemy_6_x <= writedata[9:0];
         6'h21 : enemy_6_y <= writedata[9:0];
         6'h22 : enemy_7_x <= writedata[9:0];
         6'h23 : enemy_7_y <= writedata[9:0];
         6'h24 : enemy_8_x <= writedata[9:0];
         6'h25 : enemy_8_y <= writedata[9:0];
         6'h26 : bullet_x <= writedata[9:0];
         6'h27 : bullet_y <= writedata[9:0];
         6'h28 : explosion_x <= writedata[9:0];
         6'h29 : explosion_y <= writedata[9:0];
         6'h30 : score_digit_1 <= writedata[9:0];
         6'h31 : score_digit_2 <= writedata[9:0];
         6'h32 : score_digit_3 <= writedata[9:0];
         6'h33 : score_digit_4 <= writedata[9:0];
         6'h34 : score_digit_5 <= writedata[9:0];
         6'h35 : isMusic <= writedata[0];
         6'h36 : whichClip <= writedata[1:0];
       endcase
   always_comb begin
      if (plane_y[0]) begin
	      if((hcount[10:1] - plane_x < 16) && (hcount[10:1] - plane_x > 16) && (vcount - plane_y < 16) && (vcount - plane_y[9:1] > 16)) begin // check plane sprite
	  
	      end
      end
      if (enemy_1_y[0]) begin
	      else if((hcount[10:1] - enemy_1_x < 16) && (hcount[10:1] - enemy_1_x > 16) && (vcount - enemy_1_y < 16) && (vcount - enemy_1_y[9:1] > 16)) begin // check enemy 1

	      end
      end
      if (enemy_2_y[0]) begin
	      else if((hcount[10:1] - enemy_2_x < 16) && (hcount[10:1] - enemy_2_x > 16) && (vcount - enemy_2_y < 16) && (vcount - enemy_2_y[9:1] > 16)) begin // check enemy 2

	      end
      end
      if(enemy_3_y[0]) begin
	      else if((hcount[10:1] - enemy_3_x < 16) && (hcount[10:1] - enemy_3_x > 16) && (vcount - enemy_3_y < 16) && (vcount - enemy_3_y[9:1] > 16)) begin // check enemy 3

	      end
      end
      if(enemy_4_y[0]) begin
	      else if((hcount[10:1] - enemy_4_x < 16) && (hcount[10:1] - enemy_4_x > 16) && (vcount - enemy_4_y < 16) && (vcount - enemy_4_y[9:1] > 16)) begin // check enemy 4

	      end
      end
      if(enemy_5_y[0]) begin
	      else if((hcount[10:1] - enemy_5_x < 16) && (hcount[10:1] - enemy_5_x > 16) && (vcount - enemy_5_y < 16) && (vcount - enemy_5_y[9:1] > 16)) begin // check enemy 5

	      end
      end
      if(enemy_6_y[0]) begin
	      else if((hcount[10:1] - enemy_6_x < 16) && (hcount[10:1] - enemy_6_x > 16) && (vcount - enemy_6_y < 16) && (vcount - enemy_6_y[9:1] > 16)) begin // check enemy 6

	      end
      end
      if(enemy_7_y[0]) begin
	      else if((hcount[10:1] - enemy_7_x < 16) && (hcount[10:1] - enemy_7_x > 16) && (vcount - enemy_7_y < 16) && (vcount - enemy_7_y[9:1] > 16)) begin // check enemy 7

	      end
      end
      if(enemy_8_y[0]) begin
	      else if((hcount[10:1] - enemy_8_x < 16) && (hcount[10:1] - enemy_8_x > 16) && (vcount - enemy_8_y < 16) && (vcount - enemy_8_y[9:1] > 16)) begin // check enemy 8

	      end
      end

      else if (boundary_3 == 0 && boundary_4 == 0) begin
         if  (hcount < boundary1) begin
            {VGA_R, VGA_G, VGA_B} = {8'000, 8'h00, 8'000}; // green
	 end if
         else if (hcount < boundary 2) begin
            {VGA_R, VGA_G, VGA_B} = {8'000, 8'000, 8'h00}; // blue
         end
	 else begin
	    {VGA_R, VGA_G, VGA_B} = {8'000, 8'000, 8'h00}; // green
	 end if
      end
      else begin
         if  (hcount < boundary1) begin
            {VGA_R, VGA_G, VGA_B} = {8'000, 8'h00, 8'000}; // green
	 end if
         else if (hcount < boundary2) begin
            {VGA_R, VGA_G, VGA_B} = {8'000, 8'000, 8'h00}; // blue
	 end if
         else if (hcount < boundary3) begin
            {VGA_R, VGA_G, VGA_B} = {8'000, 8'h00, 8'000}; // green
	 end if
         else if (hcount < boundary4) begin
            {VGA_R, VGA_G, VGA_B} = {8'000, 8'000, 8'h00}; // blue
	 end if
	 else begin
	    {VGA_R, VGA_G, VGA_B} = {8'000, 8'000, 8'h00}; // green
	 end if
      end if

   end
	       
endmodule

module vga_counters(
 input logic 	     clk50, reset,
 output logic [10:0] hcount,  // hcount[10:1] is pixel column
 output logic [9:0]  vcount,  // vcount[9:0] is pixel row
 output logic 	     VGA_CLK, VGA_HS, VGA_VS, VGA_BLANK_n, VGA_SYNC_n);

/*
 * 640 X 480 VGA timing for a 50 MHz clock: one pixel every other cycle
 * 
 * HCOUNT 1599 0             1279       1599 0
 *             _______________              ________
 * ___________|    Video      |____________|  Video
 * 
 * 
 * |SYNC| BP |<-- HACTIVE -->|FP|SYNC| BP |<-- HACTIVE
 *       _______________________      _____________
 * |____|       VGA_HS          |____|
 */
   // Parameters for hcount
   parameter HACTIVE      = 11'd 1280,
             HFRONT_PORCH = 11'd 32,
             HSYNC        = 11'd 192,
             HBACK_PORCH  = 11'd 96,   
             HTOTAL       = HACTIVE + HFRONT_PORCH + HSYNC +
                            HBACK_PORCH; // 1600
   
   // Parameters for vcount
   parameter VACTIVE      = 10'd 480,
             VFRONT_PORCH = 10'd 10,
             VSYNC        = 10'd 2,
             VBACK_PORCH  = 10'd 33,
             VTOTAL       = VACTIVE + VFRONT_PORCH + VSYNC +
                            VBACK_PORCH; // 525

   logic endOfLine;
   
   always_ff @(posedge clk50 or posedge reset)
     if (reset)          hcount <= 0;
     else if (endOfLine) hcount <= 0;
     else  	         hcount <= hcount + 11'd 1;

   assign endOfLine = hcount == HTOTAL - 1;
       
   logic endOfField;
   
   always_ff @(posedge clk50 or posedge reset)
     if (reset)          vcount <= 0;
     else if (endOfLine)
       if (endOfField)   vcount <= 0;
       else              vcount <= vcount + 10'd 1;

   assign endOfField = vcount == VTOTAL - 1;

   // Horizontal sync: from 0x520 to 0x5DF (0x57F)
   // 101 0010 0000 to 101 1101 1111
   assign VGA_HS = !( (hcount[10:8] == 3'b101) &
		      !(hcount[7:5] == 3'b111));
   assign VGA_VS = !( vcount[9:1] == (VACTIVE + VFRONT_PORCH) / 2);

   assign VGA_SYNC_n = 1'b0; // For putting sync on the green signal; unused
   
   // Horizontal active: 0 to 1279     Vertical active: 0 to 479
   // 101 0000 0000  1280	       01 1110 0000  480
   // 110 0011 1111  1599	       10 0000 1100  524
   assign VGA_BLANK_n = !( hcount[10] & (hcount[9] | hcount[8]) ) &
			!( vcount[9] | (vcount[8:5] == 4'b1111) );

   /* VGA_CLK is 25 MHz
    *             __    __    __
    * clk50    __|  |__|  |__|
    *        
    *             _____       __
    * hcount[0]__|     |_____|
    */
   assign VGA_CLK = hcount[0]; // 25 MHz clock: rising edge sensitive
   
endmodule
